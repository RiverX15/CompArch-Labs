module or32bit(output [31:0] out, input [31:0] in1, input [31:0] in2);
    assign out=in1|in2;
endmodule